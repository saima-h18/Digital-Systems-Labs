library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity g14_lab2 is
port(	x			: in std_logic_vector (9 downto 0);	
		y			: in std_logic_vector (9 downto 0);
		N			: in std_logic_vector (9 downto 0);
		clk		: in std_logic;
		rst		: in std_logic;
		mac		: out std_logic_vector (21 downto 0);
		ready		: out std_logic;
		counter		: out integer range 0 to 1000);
end g14_lab2;

architecture archlab2 of g14_lab2 is

signal maccounter: signed(21 downto 0);
signal count: integer range 0 to 1000 := 0;

	begin

		process(clk,rst)
		begin	
		
		if rising_edge(clk) then
			if rst = '1' then 
				maccounter <= (to_signed(0,22));
				ready <= '0';
				count <= 0;
			else
				
					maccounter <= maccounter + (signed(x) * signed(y));
					count <= count + 1;
					ready <= '0';
					
				if (count = to_integer(unsigned(N))-1) then
					ready <= '1';
				end if;				
			end if;
	
		end if;		
	end process;
	mac <= std_logic_vector(maccounter);
			counter <= count;	
end archlab2;
